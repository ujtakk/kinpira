`ifndef _NINJIN_VH_
`define _NINJIN_VH_

parameter PORT            = 32;
parameter DWIDTH          = 16;
parameter LWIDTH          = 10;
parameter IMGSIZE         = 12;

`endif
