`ifndef _RENKON_VH_
`define _RENKON_VH_

parameter RENKON_CORE    = 8;
parameter RENKON_CORELOG = 3;
parameter RENKON_NETSIZE = 11;
parameter FACCUM  = 10;
parameter BUFSIZE = 5;
parameter OUTSIZE = 8;

`endif
