
parameter DWIDTH  = 16;
parameter LWIDTH  = 10;
parameter STEP    = 10;
parameter CORE    = 8;
parameter CORELOG = 3;
parameter FACCUM  = 10;
parameter BUFSIZE = 5;
parameter IMGSIZE = 15;
parameter NETSIZE = 11;
parameter OUTSIZE = 8;
parameter N_IN    = 1;
parameter N_F1    = 16;
parameter N_F2    = 32;
parameter FSIZE   = 5;
parameter PSIZE   = 2;
