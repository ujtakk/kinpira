// % weight = "/Users/pitchw0w/work/1.hw/bhewtek/data/mnist/lenet"

`timescale 1ns/1ps

module test_gobou();
`include "gobou.vh"

  /*AUTOREGINPUT*/
  // Beginning of automatic reg inputs (for undeclared instantiated-module inputs)
  reg			clk;			// To dut0 of gobou.v
  reg			img_we;			// To dut0 of gobou.v
  reg [IMGSIZE-1:0]	input_addr;		// To dut0 of gobou.v
  reg [NETSIZE-1:0]	net_addr;		// To dut0 of gobou.v
  reg [CORELOG:0]	net_we;			// To dut0 of gobou.v
  reg [IMGSIZE-1:0]	output_addr;		// To dut0 of gobou.v
  reg signed [DWIDTH-1:0] read_img;		// To dut0 of gobou.v
  reg			req;			// To dut0 of gobou.v
  reg [LWIDTH-1:0]	total_in;		// To dut0 of gobou.v
  reg [LWIDTH-1:0]	total_out;		// To dut0 of gobou.v
  reg signed [DWIDTH-1:0] write_img;		// To dut0 of gobou.v
  reg signed [DWIDTH-1:0] write_net;		// To dut0 of gobou.v
  reg			xrst;			// To dut0 of gobou.v
  // End of automatics
  reg [DWIDTH-1:0] mem_i [2**IMGSIZE-1:0];

  /*AUTOWIRE*/
  // Beginning of automatic wires (for undeclared instantiated-module outputs)
  wire			ack;			// From dut0 of gobou.v
  wire [IMGSIZE-1:0]	mem_img_addr;		// From dut0 of gobou.v
  wire			mem_img_we;		// From dut0 of gobou.v
  wire signed [DWIDTH-1:0] write_mem_img;	// From dut0 of gobou.v
  // End of automatics
  reg [DWIDTH-1:0] mem_n0 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n1 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n2 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n3 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n4 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n5 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n6 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n7 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n8 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n9 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n10 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n11 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n12 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n13 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n14 [2**NETSIZE-1:0];
  reg [DWIDTH-1:0] mem_n15 [2**NETSIZE-1:0];

  //clock
  always
  begin
    clk = 0;
    #(STEP/2);
    clk = 1;
    #(STEP/2);
  end

  //flow
  integer i;
  initial
  begin
    xrst = 0;
    #(STEP);

    xrst = 1;
    req = 0;
    img_we = 0;
    input_addr = 0;
    output_addr = 0;
    write_img = 0;
    net_we = 0;
    net_addr = 0;
    write_net = 0;
    total_out = 0;
    total_in = 0;
    #(STEP);

    total_out = 500;
    total_in = 800;
    input_addr = 0;
    output_addr = 1000;
    read_input;
    read_weight;
    #(STEP);

    req = 1;
    #(STEP);
    req = 0;

    while(!ack) #(STEP);
    #(STEP*10);
    write_output;
    $finish();
  end

  gobou dut0(/*AUTOINST*/
	     // Outputs
	     .ack			(ack),
	     .mem_img_we		(mem_img_we),
	     .mem_img_addr		(mem_img_addr[IMGSIZE-1:0]),
	     .write_mem_img		(write_mem_img[DWIDTH-1:0]),
	     // Inputs
	     .clk			(clk),
	     .xrst			(xrst),
	     .req			(req),
	     .img_we			(img_we),
	     .input_addr		(input_addr[IMGSIZE-1:0]),
	     .output_addr		(output_addr[IMGSIZE-1:0]),
	     .write_img			(write_img[DWIDTH-1:0]),
	     .net_we			(net_we[CORELOG:0]),
	     .net_addr			(net_addr[NETSIZE-1:0]),
	     .write_net			(write_net[DWIDTH-1:0]),
	     .total_out			(total_out[LWIDTH-1:0]),
	     .total_in			(total_in[LWIDTH-1:0]),
	     .read_img			(read_img[DWIDTH-1:0]));

  task read_input;
    begin // {{{
      $readmemh(
        "test_gobou_input.dat",
        mem_i,
        0,
        799
      );
      img_we = 1;
        #(STEP);
      for (i=0; i<2**IMGSIZE; i=i+1)
      begin
        input_addr = i;
        #(STEP);
        write_img = mem_i[i];
        #(STEP);
      end
      #(STEP);
      img_we = 0;
      input_addr = 0;
      write_img = 0;
    end // }}}
  endtask

  task read_input_direct;
    begin // {{{
      $readmemh(
        "test_gobou_input.dat",
        dut0.mem_img.mem,
        0,
        799
      );
    end // }}}
  endtask

  task read_weight;
    begin // {{{
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data0.bin",
        mem_n0,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data1.bin",
        mem_n1,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data2.bin",
        mem_n2,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data3.bin",
        mem_n3,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data4.bin",
        mem_n4,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data5.bin",
        mem_n5,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data6.bin",
        mem_n6,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data7.bin",
        mem_n7,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data8.bin",
        mem_n8,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data9.bin",
        mem_n9,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data10.bin",
        mem_n10,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data11.bin",
        mem_n11,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data12.bin",
        mem_n12,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data13.bin",
        mem_n13,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data14.bin",
        mem_n14,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data15.bin",
        mem_n15,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data16.bin",
        mem_n0,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data17.bin",
        mem_n1,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data18.bin",
        mem_n2,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data19.bin",
        mem_n3,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data20.bin",
        mem_n4,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data21.bin",
        mem_n5,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data22.bin",
        mem_n6,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data23.bin",
        mem_n7,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data24.bin",
        mem_n8,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data25.bin",
        mem_n9,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data26.bin",
        mem_n10,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data27.bin",
        mem_n11,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data28.bin",
        mem_n12,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data29.bin",
        mem_n13,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data30.bin",
        mem_n14,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data31.bin",
        mem_n15,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data32.bin",
        mem_n0,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data33.bin",
        mem_n1,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data34.bin",
        mem_n2,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data35.bin",
        mem_n3,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data36.bin",
        mem_n4,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data37.bin",
        mem_n5,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data38.bin",
        mem_n6,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data39.bin",
        mem_n7,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data40.bin",
        mem_n8,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data41.bin",
        mem_n9,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data42.bin",
        mem_n10,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data43.bin",
        mem_n11,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data44.bin",
        mem_n12,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data45.bin",
        mem_n13,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data46.bin",
        mem_n14,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data47.bin",
        mem_n15,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data48.bin",
        mem_n0,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data49.bin",
        mem_n1,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data50.bin",
        mem_n2,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data51.bin",
        mem_n3,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data52.bin",
        mem_n4,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data53.bin",
        mem_n5,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data54.bin",
        mem_n6,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data55.bin",
        mem_n7,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data56.bin",
        mem_n8,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data57.bin",
        mem_n9,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data58.bin",
        mem_n10,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data59.bin",
        mem_n11,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data60.bin",
        mem_n12,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data61.bin",
        mem_n13,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data62.bin",
        mem_n14,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data63.bin",
        mem_n15,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data64.bin",
        mem_n0,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data65.bin",
        mem_n1,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data66.bin",
        mem_n2,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data67.bin",
        mem_n3,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data68.bin",
        mem_n4,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data69.bin",
        mem_n5,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data70.bin",
        mem_n6,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data71.bin",
        mem_n7,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data72.bin",
        mem_n8,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data73.bin",
        mem_n9,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data74.bin",
        mem_n10,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data75.bin",
        mem_n11,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data76.bin",
        mem_n12,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data77.bin",
        mem_n13,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data78.bin",
        mem_n14,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data79.bin",
        mem_n15,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data80.bin",
        mem_n0,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data81.bin",
        mem_n1,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data82.bin",
        mem_n2,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data83.bin",
        mem_n3,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data84.bin",
        mem_n4,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data85.bin",
        mem_n5,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data86.bin",
        mem_n6,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data87.bin",
        mem_n7,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data88.bin",
        mem_n8,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data89.bin",
        mem_n9,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data90.bin",
        mem_n10,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data91.bin",
        mem_n11,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data92.bin",
        mem_n12,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data93.bin",
        mem_n13,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data94.bin",
        mem_n14,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data95.bin",
        mem_n15,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data96.bin",
        mem_n0,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data97.bin",
        mem_n1,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data98.bin",
        mem_n2,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data99.bin",
        mem_n3,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data100.bin",
        mem_n4,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data101.bin",
        mem_n5,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data102.bin",
        mem_n6,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data103.bin",
        mem_n7,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data104.bin",
        mem_n8,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data105.bin",
        mem_n9,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data106.bin",
        mem_n10,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data107.bin",
        mem_n11,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data108.bin",
        mem_n12,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data109.bin",
        mem_n13,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data110.bin",
        mem_n14,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data111.bin",
        mem_n15,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data112.bin",
        mem_n0,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data113.bin",
        mem_n1,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data114.bin",
        mem_n2,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data115.bin",
        mem_n3,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data116.bin",
        mem_n4,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data117.bin",
        mem_n5,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data118.bin",
        mem_n6,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data119.bin",
        mem_n7,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data120.bin",
        mem_n8,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data121.bin",
        mem_n9,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data122.bin",
        mem_n10,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data123.bin",
        mem_n11,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data124.bin",
        mem_n12,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data125.bin",
        mem_n13,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data126.bin",
        mem_n14,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data127.bin",
        mem_n15,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data128.bin",
        mem_n0,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data129.bin",
        mem_n1,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data130.bin",
        mem_n2,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data131.bin",
        mem_n3,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data132.bin",
        mem_n4,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data133.bin",
        mem_n5,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data134.bin",
        mem_n6,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data135.bin",
        mem_n7,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data136.bin",
        mem_n8,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data137.bin",
        mem_n9,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data138.bin",
        mem_n10,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data139.bin",
        mem_n11,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data140.bin",
        mem_n12,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data141.bin",
        mem_n13,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data142.bin",
        mem_n14,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data143.bin",
        mem_n15,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data144.bin",
        mem_n0,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data145.bin",
        mem_n1,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data146.bin",
        mem_n2,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data147.bin",
        mem_n3,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data148.bin",
        mem_n4,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data149.bin",
        mem_n5,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data150.bin",
        mem_n6,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data151.bin",
        mem_n7,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data152.bin",
        mem_n8,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data153.bin",
        mem_n9,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data154.bin",
        mem_n10,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data155.bin",
        mem_n11,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data156.bin",
        mem_n12,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data157.bin",
        mem_n13,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data158.bin",
        mem_n14,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data159.bin",
        mem_n15,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data160.bin",
        mem_n0,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data161.bin",
        mem_n1,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data162.bin",
        mem_n2,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data163.bin",
        mem_n3,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data164.bin",
        mem_n4,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data165.bin",
        mem_n5,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data166.bin",
        mem_n6,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data167.bin",
        mem_n7,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data168.bin",
        mem_n8,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data169.bin",
        mem_n9,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data170.bin",
        mem_n10,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data171.bin",
        mem_n11,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data172.bin",
        mem_n12,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data173.bin",
        mem_n13,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data174.bin",
        mem_n14,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data175.bin",
        mem_n15,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data176.bin",
        mem_n0,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data177.bin",
        mem_n1,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data178.bin",
        mem_n2,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data179.bin",
        mem_n3,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data180.bin",
        mem_n4,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data181.bin",
        mem_n5,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data182.bin",
        mem_n6,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data183.bin",
        mem_n7,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data184.bin",
        mem_n8,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data185.bin",
        mem_n9,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data186.bin",
        mem_n10,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data187.bin",
        mem_n11,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data188.bin",
        mem_n12,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data189.bin",
        mem_n13,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data190.bin",
        mem_n14,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data191.bin",
        mem_n15,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data192.bin",
        mem_n0,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data193.bin",
        mem_n1,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data194.bin",
        mem_n2,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data195.bin",
        mem_n3,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data196.bin",
        mem_n4,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data197.bin",
        mem_n5,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data198.bin",
        mem_n6,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data199.bin",
        mem_n7,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data200.bin",
        mem_n8,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data201.bin",
        mem_n9,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data202.bin",
        mem_n10,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data203.bin",
        mem_n11,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data204.bin",
        mem_n12,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data205.bin",
        mem_n13,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data206.bin",
        mem_n14,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data207.bin",
        mem_n15,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data208.bin",
        mem_n0,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data209.bin",
        mem_n1,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data210.bin",
        mem_n2,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data211.bin",
        mem_n3,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data212.bin",
        mem_n4,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data213.bin",
        mem_n5,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data214.bin",
        mem_n6,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data215.bin",
        mem_n7,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data216.bin",
        mem_n8,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data217.bin",
        mem_n9,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data218.bin",
        mem_n10,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data219.bin",
        mem_n11,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data220.bin",
        mem_n12,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data221.bin",
        mem_n13,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data222.bin",
        mem_n14,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data223.bin",
        mem_n15,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data224.bin",
        mem_n0,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data225.bin",
        mem_n1,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data226.bin",
        mem_n2,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data227.bin",
        mem_n3,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data228.bin",
        mem_n4,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data229.bin",
        mem_n5,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data230.bin",
        mem_n6,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data231.bin",
        mem_n7,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data232.bin",
        mem_n8,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data233.bin",
        mem_n9,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data234.bin",
        mem_n10,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data235.bin",
        mem_n11,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data236.bin",
        mem_n12,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data237.bin",
        mem_n13,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data238.bin",
        mem_n14,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data239.bin",
        mem_n15,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data240.bin",
        mem_n0,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data241.bin",
        mem_n1,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data242.bin",
        mem_n2,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data243.bin",
        mem_n3,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data244.bin",
        mem_n4,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data245.bin",
        mem_n5,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data246.bin",
        mem_n6,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data247.bin",
        mem_n7,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data248.bin",
        mem_n8,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data249.bin",
        mem_n9,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data250.bin",
        mem_n10,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data251.bin",
        mem_n11,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data252.bin",
        mem_n12,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data253.bin",
        mem_n13,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data254.bin",
        mem_n14,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data255.bin",
        mem_n15,
        7695,
        8207
      );

      net_we = 5'd1;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n0[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd2;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n1[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd3;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n2[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd4;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n3[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd5;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n4[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd6;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n5[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd7;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n6[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd8;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n7[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd9;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n8[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd10;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n9[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd11;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n10[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd12;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n11[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd13;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n12[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd14;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n13[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd15;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n14[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
      net_we = 5'd16;
      #(STEP);
      for (i=0; i<2**NETSIZE; i=i+1)
      begin
        net_addr = i;
        #(STEP);
        write_net = mem_n15[i];
        #(STEP);
      end
      net_we = 5'd0;
      net_addr = 0;
      write_net = 0;
    end // }}}
  endtask

  task read_weight_direct;
    begin // {{{
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data0.bin",
        dut0.mem_net0.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data1.bin",
        dut0.mem_net1.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data2.bin",
        dut0.mem_net2.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data3.bin",
        dut0.mem_net3.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data4.bin",
        dut0.mem_net4.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data5.bin",
        dut0.mem_net5.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data6.bin",
        dut0.mem_net6.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data7.bin",
        dut0.mem_net7.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data8.bin",
        dut0.mem_net8.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data9.bin",
        dut0.mem_net9.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data10.bin",
        dut0.mem_net10.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data11.bin",
        dut0.mem_net11.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data12.bin",
        dut0.mem_net12.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data13.bin",
        dut0.mem_net13.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data14.bin",
        dut0.mem_net14.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data15.bin",
        dut0.mem_net15.mem,
        0,
        512
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data16.bin",
        dut0.mem_net0.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data17.bin",
        dut0.mem_net1.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data18.bin",
        dut0.mem_net2.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data19.bin",
        dut0.mem_net3.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data20.bin",
        dut0.mem_net4.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data21.bin",
        dut0.mem_net5.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data22.bin",
        dut0.mem_net6.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data23.bin",
        dut0.mem_net7.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data24.bin",
        dut0.mem_net8.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data25.bin",
        dut0.mem_net9.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data26.bin",
        dut0.mem_net10.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data27.bin",
        dut0.mem_net11.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data28.bin",
        dut0.mem_net12.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data29.bin",
        dut0.mem_net13.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data30.bin",
        dut0.mem_net14.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data31.bin",
        dut0.mem_net15.mem,
        513,
        1025
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data32.bin",
        dut0.mem_net0.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data33.bin",
        dut0.mem_net1.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data34.bin",
        dut0.mem_net2.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data35.bin",
        dut0.mem_net3.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data36.bin",
        dut0.mem_net4.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data37.bin",
        dut0.mem_net5.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data38.bin",
        dut0.mem_net6.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data39.bin",
        dut0.mem_net7.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data40.bin",
        dut0.mem_net8.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data41.bin",
        dut0.mem_net9.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data42.bin",
        dut0.mem_net10.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data43.bin",
        dut0.mem_net11.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data44.bin",
        dut0.mem_net12.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data45.bin",
        dut0.mem_net13.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data46.bin",
        dut0.mem_net14.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data47.bin",
        dut0.mem_net15.mem,
        1026,
        1538
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data48.bin",
        dut0.mem_net0.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data49.bin",
        dut0.mem_net1.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data50.bin",
        dut0.mem_net2.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data51.bin",
        dut0.mem_net3.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data52.bin",
        dut0.mem_net4.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data53.bin",
        dut0.mem_net5.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data54.bin",
        dut0.mem_net6.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data55.bin",
        dut0.mem_net7.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data56.bin",
        dut0.mem_net8.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data57.bin",
        dut0.mem_net9.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data58.bin",
        dut0.mem_net10.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data59.bin",
        dut0.mem_net11.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data60.bin",
        dut0.mem_net12.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data61.bin",
        dut0.mem_net13.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data62.bin",
        dut0.mem_net14.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data63.bin",
        dut0.mem_net15.mem,
        1539,
        2051
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data64.bin",
        dut0.mem_net0.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data65.bin",
        dut0.mem_net1.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data66.bin",
        dut0.mem_net2.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data67.bin",
        dut0.mem_net3.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data68.bin",
        dut0.mem_net4.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data69.bin",
        dut0.mem_net5.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data70.bin",
        dut0.mem_net6.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data71.bin",
        dut0.mem_net7.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data72.bin",
        dut0.mem_net8.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data73.bin",
        dut0.mem_net9.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data74.bin",
        dut0.mem_net10.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data75.bin",
        dut0.mem_net11.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data76.bin",
        dut0.mem_net12.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data77.bin",
        dut0.mem_net13.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data78.bin",
        dut0.mem_net14.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data79.bin",
        dut0.mem_net15.mem,
        2052,
        2564
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data80.bin",
        dut0.mem_net0.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data81.bin",
        dut0.mem_net1.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data82.bin",
        dut0.mem_net2.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data83.bin",
        dut0.mem_net3.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data84.bin",
        dut0.mem_net4.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data85.bin",
        dut0.mem_net5.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data86.bin",
        dut0.mem_net6.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data87.bin",
        dut0.mem_net7.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data88.bin",
        dut0.mem_net8.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data89.bin",
        dut0.mem_net9.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data90.bin",
        dut0.mem_net10.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data91.bin",
        dut0.mem_net11.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data92.bin",
        dut0.mem_net12.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data93.bin",
        dut0.mem_net13.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data94.bin",
        dut0.mem_net14.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data95.bin",
        dut0.mem_net15.mem,
        2565,
        3077
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data96.bin",
        dut0.mem_net0.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data97.bin",
        dut0.mem_net1.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data98.bin",
        dut0.mem_net2.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data99.bin",
        dut0.mem_net3.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data100.bin",
        dut0.mem_net4.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data101.bin",
        dut0.mem_net5.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data102.bin",
        dut0.mem_net6.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data103.bin",
        dut0.mem_net7.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data104.bin",
        dut0.mem_net8.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data105.bin",
        dut0.mem_net9.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data106.bin",
        dut0.mem_net10.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data107.bin",
        dut0.mem_net11.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data108.bin",
        dut0.mem_net12.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data109.bin",
        dut0.mem_net13.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data110.bin",
        dut0.mem_net14.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data111.bin",
        dut0.mem_net15.mem,
        3078,
        3590
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data112.bin",
        dut0.mem_net0.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data113.bin",
        dut0.mem_net1.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data114.bin",
        dut0.mem_net2.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data115.bin",
        dut0.mem_net3.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data116.bin",
        dut0.mem_net4.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data117.bin",
        dut0.mem_net5.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data118.bin",
        dut0.mem_net6.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data119.bin",
        dut0.mem_net7.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data120.bin",
        dut0.mem_net8.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data121.bin",
        dut0.mem_net9.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data122.bin",
        dut0.mem_net10.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data123.bin",
        dut0.mem_net11.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data124.bin",
        dut0.mem_net12.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data125.bin",
        dut0.mem_net13.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data126.bin",
        dut0.mem_net14.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data127.bin",
        dut0.mem_net15.mem,
        3591,
        4103
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data128.bin",
        dut0.mem_net0.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data129.bin",
        dut0.mem_net1.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data130.bin",
        dut0.mem_net2.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data131.bin",
        dut0.mem_net3.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data132.bin",
        dut0.mem_net4.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data133.bin",
        dut0.mem_net5.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data134.bin",
        dut0.mem_net6.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data135.bin",
        dut0.mem_net7.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data136.bin",
        dut0.mem_net8.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data137.bin",
        dut0.mem_net9.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data138.bin",
        dut0.mem_net10.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data139.bin",
        dut0.mem_net11.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data140.bin",
        dut0.mem_net12.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data141.bin",
        dut0.mem_net13.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data142.bin",
        dut0.mem_net14.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data143.bin",
        dut0.mem_net15.mem,
        4104,
        4616
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data144.bin",
        dut0.mem_net0.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data145.bin",
        dut0.mem_net1.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data146.bin",
        dut0.mem_net2.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data147.bin",
        dut0.mem_net3.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data148.bin",
        dut0.mem_net4.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data149.bin",
        dut0.mem_net5.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data150.bin",
        dut0.mem_net6.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data151.bin",
        dut0.mem_net7.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data152.bin",
        dut0.mem_net8.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data153.bin",
        dut0.mem_net9.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data154.bin",
        dut0.mem_net10.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data155.bin",
        dut0.mem_net11.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data156.bin",
        dut0.mem_net12.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data157.bin",
        dut0.mem_net13.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data158.bin",
        dut0.mem_net14.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data159.bin",
        dut0.mem_net15.mem,
        4617,
        5129
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data160.bin",
        dut0.mem_net0.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data161.bin",
        dut0.mem_net1.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data162.bin",
        dut0.mem_net2.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data163.bin",
        dut0.mem_net3.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data164.bin",
        dut0.mem_net4.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data165.bin",
        dut0.mem_net5.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data166.bin",
        dut0.mem_net6.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data167.bin",
        dut0.mem_net7.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data168.bin",
        dut0.mem_net8.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data169.bin",
        dut0.mem_net9.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data170.bin",
        dut0.mem_net10.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data171.bin",
        dut0.mem_net11.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data172.bin",
        dut0.mem_net12.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data173.bin",
        dut0.mem_net13.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data174.bin",
        dut0.mem_net14.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data175.bin",
        dut0.mem_net15.mem,
        5130,
        5642
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data176.bin",
        dut0.mem_net0.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data177.bin",
        dut0.mem_net1.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data178.bin",
        dut0.mem_net2.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data179.bin",
        dut0.mem_net3.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data180.bin",
        dut0.mem_net4.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data181.bin",
        dut0.mem_net5.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data182.bin",
        dut0.mem_net6.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data183.bin",
        dut0.mem_net7.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data184.bin",
        dut0.mem_net8.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data185.bin",
        dut0.mem_net9.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data186.bin",
        dut0.mem_net10.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data187.bin",
        dut0.mem_net11.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data188.bin",
        dut0.mem_net12.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data189.bin",
        dut0.mem_net13.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data190.bin",
        dut0.mem_net14.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data191.bin",
        dut0.mem_net15.mem,
        5643,
        6155
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data192.bin",
        dut0.mem_net0.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data193.bin",
        dut0.mem_net1.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data194.bin",
        dut0.mem_net2.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data195.bin",
        dut0.mem_net3.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data196.bin",
        dut0.mem_net4.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data197.bin",
        dut0.mem_net5.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data198.bin",
        dut0.mem_net6.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data199.bin",
        dut0.mem_net7.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data200.bin",
        dut0.mem_net8.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data201.bin",
        dut0.mem_net9.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data202.bin",
        dut0.mem_net10.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data203.bin",
        dut0.mem_net11.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data204.bin",
        dut0.mem_net12.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data205.bin",
        dut0.mem_net13.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data206.bin",
        dut0.mem_net14.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data207.bin",
        dut0.mem_net15.mem,
        6156,
        6668
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data208.bin",
        dut0.mem_net0.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data209.bin",
        dut0.mem_net1.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data210.bin",
        dut0.mem_net2.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data211.bin",
        dut0.mem_net3.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data212.bin",
        dut0.mem_net4.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data213.bin",
        dut0.mem_net5.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data214.bin",
        dut0.mem_net6.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data215.bin",
        dut0.mem_net7.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data216.bin",
        dut0.mem_net8.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data217.bin",
        dut0.mem_net9.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data218.bin",
        dut0.mem_net10.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data219.bin",
        dut0.mem_net11.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data220.bin",
        dut0.mem_net12.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data221.bin",
        dut0.mem_net13.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data222.bin",
        dut0.mem_net14.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data223.bin",
        dut0.mem_net15.mem,
        6669,
        7181
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data224.bin",
        dut0.mem_net0.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data225.bin",
        dut0.mem_net1.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data226.bin",
        dut0.mem_net2.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data227.bin",
        dut0.mem_net3.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data228.bin",
        dut0.mem_net4.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data229.bin",
        dut0.mem_net5.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data230.bin",
        dut0.mem_net6.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data231.bin",
        dut0.mem_net7.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data232.bin",
        dut0.mem_net8.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data233.bin",
        dut0.mem_net9.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data234.bin",
        dut0.mem_net10.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data235.bin",
        dut0.mem_net11.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data236.bin",
        dut0.mem_net12.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data237.bin",
        dut0.mem_net13.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data238.bin",
        dut0.mem_net14.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data239.bin",
        dut0.mem_net15.mem,
        7182,
        7694
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data240.bin",
        dut0.mem_net0.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data241.bin",
        dut0.mem_net1.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data242.bin",
        dut0.mem_net2.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data243.bin",
        dut0.mem_net3.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data244.bin",
        dut0.mem_net4.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data245.bin",
        dut0.mem_net5.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data246.bin",
        dut0.mem_net6.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data247.bin",
        dut0.mem_net7.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data248.bin",
        dut0.mem_net8.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data249.bin",
        dut0.mem_net9.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data250.bin",
        dut0.mem_net10.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data251.bin",
        dut0.mem_net11.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data252.bin",
        dut0.mem_net12.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data253.bin",
        dut0.mem_net13.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data254.bin",
        dut0.mem_net14.mem,
        7695,
        8207
      );
      $readmemb(
        "/home/work/takau/bhewtek/data/mnist/lenet/bwb_3/data255.bin",
        dut0.mem_net15.mem,
        7695,
        8207
      );
    end // }}}
  endtask

  task write_output;
    integer fd;
    integer i;
    integer out_size;
    begin // {{{
      fd = $fopen("test_gobou.dat", "w");
      out_size = 500;
      for (i=1000; i<1000+out_size; i=i+1)
        $fdisplay(fd, "%0d", dut0.mem_img.mem[i]);
      $fclose(fd);
    end // }}}
  endtask

  //display
  always
  begin
    #(STEP/2-1);
    $display(
      "%5d: ", $time/STEP,
      "%d ", dut0.ctrl.ctrl_core.r_state,
      "| ",
      "%d ", clk,
      "%d ", xrst,
      "%d ", req,
      "%d ", img_we,
      "%3d ", input_addr,
      "%3d ", output_addr,
      "%d ", write_img,
      "%d ", net_we,
      "%3d ", net_addr,
      "%3d ", write_net,
      "%3d ", total_out,
      "%3d ", total_in,
      "| ",
      "%d ", ack,
      "%d ", read_img,
      "| ",
      "%d ", dut0.ctrl.out_core_valid,
      "%d ", dut0.ctrl.out_mac_valid,
      "%d ", dut0.ctrl.out_bias_valid,
      "%d ", dut0.ctrl.out_relu_valid,
      ": ",
      "%d ", dut0.core0.mac_oe,
      "%d ", dut0.core0.bias_oe,
      "%d ", dut0.core0.relu_oe,
      "%d ", dut0.serial_we,
      "| ",
      "%d ", dut0.mem_img_we,
      "%4d ", dut0.mem_img_addr,
      "%3d ", dut0.write_mem_img,
      "%3d ", dut0.write_result,
      "%d ", dut0.mem_img.mem[1000],
      "| ",
      "%d ", dut0.core0.accum_we,
      "%x ", dut0.core0.pixel,
      "%d ", dut0.core0.weight,
      "%d ", dut0.core0.bias.r_bias,
      "%d ", dut0.core0.dotted,
      "%d ", dut0.core0.biased,
      "%d ", dut0.core0.result,
      "%d ", dut0.serial.r_data0,
      "|"
    );
    #(STEP/2+1);
  end

endmodule
