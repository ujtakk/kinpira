`ifndef _GOBOU_VH_
`define _GOBOU_VH_

parameter GOBOU_CORE    = 16;
parameter GOBOU_CORELOG = 4;
parameter GOBOU_NETSIZE = 14;

`endif
